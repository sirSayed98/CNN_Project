-- 
-- Layer counter
-- Depth counter
-- Filter counter 