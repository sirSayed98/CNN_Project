
library ieee;
use ieee.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity system is
	port(
		clk : in std_logic
	    );
end entity system;

ARCHITECTURE system_arch OF system is

end system_arch;